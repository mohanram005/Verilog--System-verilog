//gate level using gate with instatation
module gate(input a,b,
            output c);
  and a1(c,a,b);
  
endmodule
