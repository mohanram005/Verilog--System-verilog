interface operation;
  
  logic d;
  logic clk;
  logic reset;
  bit q;
  
endinterface
