interface operation;
  
  logic x,y,z;
  logic sum,carry;
  
endinterface
  
