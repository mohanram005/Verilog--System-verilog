class transaction;
  
  rand logic d;
  rand bit clk;
  rand bit reset;
  bit q;
  
endclass
