
/data flow level using continous assignment
module gate(input a,b,
            output c);
  assign c = a & b;
  
endmodule
