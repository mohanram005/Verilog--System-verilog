class transaction;
rand logic x;
rand logic y;
rand logic z;

bit sum;
bit carry;
  
endclass
